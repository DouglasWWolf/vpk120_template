//================================================================================================
// Version  Date         Who  What
// -----------------------------------------------------------------------------------------------
//   1.0.0  18-Aug-25    DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0; 
localparam RTL_TYPE      = 81825;
localparam RTL_SUBTYPE   = 0;

